module NPC (
    input  clk,
    input  reset
);
endmodule
