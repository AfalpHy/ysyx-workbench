import "DPI-C" function void set_skip_ref_inst();
import "DPI-C" function void lsu_record0(
  int addr,
  int data,
  int delay
);
import "DPI-C" function void lsu_record1(
  int addr,
  int data,
  int mask,
  int delay
);
module ysyx_25010008_LSU (
    input clock,
    input reset,

    input suffix_b,
    input suffix_h,
    input sext,

    input ren,
    input wen,

    input [31:0] addr,
    input [31:0] wsrc,
    input [31:0] exu_r_wdata,
    output reg [31:0] r_wdata,
    output reg block,

    output reg arvalid,
    output [31:0] araddr,
    output [2:0] arsize,
    input arready,

    output reg rready,
    input [31:0] rdata,
    input [1:0] rresp,
    input rvalid,

    output reg awvalid,
    output [31:0] awaddr,
    output [2:0] awsize,
    input awready,

    output reg wvalid,
    output [31:0] wdata,
    output [3:0] wstrb,
    input wready,

    output reg bready,
    input [1:0] bresp,
    input bvalid
);

  reg [31:0] addr_q;
  reg suffix_b_q;
  reg suffix_h_q;
  reg sext_q;

  assign araddr = addr_q;
  assign arsize = suffix_b_q ? 0 : suffix_h_q ? 1 : 2;

  assign awaddr = addr_q;
  assign awsize = suffix_b_q ? 0 : suffix_h_q ? 1 : 2;

  assign wdata  = (suffix_b_q | suffix_h_q) ? (wsrc << {addr_q[1:0], 3'b0}) : wsrc;
  assign wstrb  = (suffix_b_q ? 4'b0001 : (suffix_h_q ? 4'b0011 : 4'b1111)) << addr_q[1:0];

  wire [31:0] real_rdata = (suffix_b_q | suffix_h_q) ? (rdata >> {addr_q[1:0], 3'b0}) : rdata;
  wire [31:0] sextb = {{24{real_rdata[7]}}, real_rdata[7:0]};
  wire [31:0] sexth = {{16{real_rdata[15]}}, real_rdata[15:0]};
  wire [31:0] sign_data = suffix_b_q ? sextb : sexth;
  wire [31:0] extb = {24'b0, real_rdata[7:0]};
  wire [31:0] exth = {16'b0, real_rdata[15:0]};
  wire [31:0] unsign_data = suffix_b_q ? extb : (suffix_h_q ? exth : real_rdata);

  integer delay;

  always @(posedge clock) begin
    if (reset) begin
      arvalid <= 0;
      rready  <= 0;

      awvalid <= 0;
      wvalid  <= 0;
      bready  <= 0;

      block   <= 0;
      delay = 0;
    end else begin
      if (block) begin
        delay = delay + 1;

        if (arvalid & arready) begin
          if (araddr[31:12] == 20'h1_0000 || araddr[31:24] == 8'h02 || araddr[31:12] == 20'h1_0001 || araddr[31:12] == 20'h1_0002 || araddr[31:12] == 20'h1_0011)
            set_skip_ref_inst();  //uart clint spi gpio ps2
          rready  <= 1;
          arvalid <= 0;
        end

        if (rready & rvalid) begin
          rready  <= 0;
          r_wdata <= sext_q ? sign_data : unsign_data;
          block   <= 0;
          lsu_record0(araddr, sext_q ? sign_data : unsign_data, delay);
          delay = 0;
        end

        if (awvalid & awready) begin
          if (awaddr[31:12] == 20'h1_0000 || araddr[31:12] == 20'h1_0001 || araddr[31:12] == 20'h1_0002 || araddr[31:24] == 8'h21)
            set_skip_ref_inst();  //uart spi gpio vga
          awvalid <= 0;
        end

        if (wvalid & wready) begin
          wvalid <= 0;
          bready <= 1;
        end

        if (bready & bvalid) begin
          bready <= 0;
          block  <= 0;
          lsu_record1(araddr, wdata, {28'b0, wstrb}, delay);
          delay = 0;
        end
      end else begin
        if (ren | wen) begin
          block <= 1;
          addr_q <= addr;
          suffix_b_q <= suffix_b;
          suffix_h_q <= suffix_h;
          sext_q <= sext;
        end

        r_wdata <= exu_r_wdata;

        if (ren) begin
          arvalid <= 1;
        end

        if (wen) begin
          // must assert in the same time for sdram axi
          awvalid <= 1;
          wvalid  <= 1;
        end
      end
    end
  end

endmodule
